module foobari (input integer a, input integer b, output integer c);
 assign c =  a*b;	
endmodule : foobari